library verilog;
use verilog.vl_types.all;
entity Lab2_tb is
end Lab2_tb;
