library verilog;
use verilog.vl_types.all;
entity sub_tb is
end sub_tb;
