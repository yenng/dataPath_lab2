library verilog;
use verilog.vl_types.all;
entity instructionSetOperation_tb is
end instructionSetOperation_tb;
