library verilog;
use verilog.vl_types.all;
entity dataPath_tb is
end dataPath_tb;
