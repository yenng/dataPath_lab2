module dataPath(
	input IRload,JMPmux, PCload, Meminst, MemWr, Aload, Reset, Clock, Sub,In,
	input [1:0] Asel,
	input [7:0] Input,
	output Aeq0, Apos,
	output [4:0] Address,
	output wire [2:0] IR,
	output [7:0] Output, RAM_Q);
	
		
	instructionCycleOperation 	part1(IRload,JMPmux,PCload,Meminst,Clock,Reset,RAM_Q,IR,Address);
	memRAM						part2(Clock,In,Output,Address,MemWr,RAM_Q);
	instructionSetOperation		part3(Aload, Reset, Clock, Sub,Asel,Input,RAM_Q,Aeq0,Apos,Output);

endmodule 